module ysyx_24120006_EXU(

);
endmodule